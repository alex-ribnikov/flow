

#
# Copyright      : Broadcom Limited 2019
# Target process : TSMC 5nm Process
#  
#
# Description    : 17M w/ 1-M1 1-Mx 1-Mxb 1-Mxe 1-Mya 1-Myb 5-My 2-Myy 2-Myx 2-Mr plus UTRDL
# Tracking       : Enterprise
#  

VERSION 5.8 ;

PROPERTYDEFINITIONS

  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA2_4X4_USER LAYER VIA2 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA3_4X4_USER LAYER VIA3 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA4_4X4_USER LAYER VIA4 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 ;" ;  
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA5_4X4_USER LAYER VIA5 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA6_4X4_USER LAYER VIA6 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA7_4X4_USER LAYER VIA7 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 2 ;" ;

  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA8_4X4_USER LAYER VIA8 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 ;" ; 
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA8_2X2_BIG_USER LAYER VIA8 CUTCLASS VSINGLECUT58 ROWCOL 2 2 XPITCH 2 YPITCH 2 ;" ; 
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA9_4X4_USER LAYER VIA9 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA10_4X4_USER LAYER VIA10 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA11_3X4_USER LAYER VIA11 CUTCLASS VSINGLECUT ROWCOL 3 4 XPITCH 3 YPITCH 2 MAXCELLEXTENSION 2 ;" ;  
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA12_3X1_USER LAYER VIA12 CUTCLASS VSINGLECUT ROWCOL 3 1 MAXXLINEEND 2 2 ;" ;    

  LIBRARY LEF58_STACKVIARULE STRING "STACKVIARULE MY_VP   VIA2_4X4_USER VIA3_4X4_USER VIA4_4X4_USER VIA5_4X4_USER VIA6_4X4_USER VIA7_4X4_USER VIA8_4X4_USER VIA9_4X4_USER VIA10_4X4_USER VIA11_3X4_USER VIA12_3X1_USER ;" ;
  
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA6_4X1_USER LAYER VIA6 CUTCLASS VSINGLECUT ROWCOL 4 1 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA7_1X4_USER LAYER VIA7 CUTCLASS VSINGLECUT ROWCOL 1 4 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 2 ;" ;  
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA8_4X1_USER LAYER VIA8 CUTCLASS VSINGLECUT ROWCOL 4 1 XPITCH 2 YPITCH 2 ;" ; 
    
  LIBRARY LEF58_STACKVIARULE STRING "STACKVIARULE MY_VP2  VIA2_4X4_USER VIA3_4X4_USER VIA4_4X4_USER VIA5_4X4_USER VIA6_4X4_USER VIA7_4X4_USER VIA8_4X1_USER ;" ;  

#  Enhance M2-M3-M4 ladder
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA2_4X8_USER LAYER VIA2 CUTCLASS VSINGLECUT ROWCOL 4 8 XPITCH 2 YPITCH 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA3_4X8_USER LAYER VIA3 CUTCLASS VSINGLECUT ROWCOL 4 8 XPITCH 2 YPITCH 2 ;" ;
#  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA4_4X4_USER LAYER VIA4 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 ;" ;  
#  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA5_4X4_USER LAYER VIA5 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 2 ;" ;

  LIBRARY LEF58_STACKVIARULE STRING "STACKVIARULE MY_VP3  VIA2_4X8_USER VIA3_4X8_USER VIA4_4X4_USER VIA5_4X4_USER VIA6_4X4_USER VIA7_4X4_USER VIA8_4X1_USER ;" ;    

  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA2_4X8_3X_USER LAYER VIA2 CUTCLASS VSINGLECUT ROWCOL 4 8 XPITCH 3 YPITCH 2 ;" ;
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA3_4X8_3X_USER LAYER VIA3 CUTCLASS VSINGLECUT ROWCOL 4 8 XPITCH 3 YPITCH 2 ;" ;
#  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA4_4X4_USER LAYER VIA4 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 ;" ;  
#  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA5_4X4_USER LAYER VIA5 CUTCLASS VSINGLECUT ROWCOL 4 4 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 2 ;" ;

  LIBRARY LEF58_STACKVIARULE STRING "STACKVIARULE MY_VP4  VIA2_4X8_3X_USER VIA3_4X8_3X_USER VIA4_4X4_USER VIA5_4X4_USER VIA6_4X4_USER VIA7_4X4_USER VIA8_4X1_USER ;" ;    
  
  # Heigher layers
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA8_4X3_USER LAYER VIA8 CUTCLASS VSINGLECUT ROWCOL 4 3 XPITCH 2 YPITCH 2 ;" ;   
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA9_3X4_USER LAYER VIA9 CUTCLASS VSINGLECUT ROWCOL 3 4 XPITCH 3 YPITCH 2 ;" ;  
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA10_3X1_USER LAYER VIA10 CUTCLASS VSINGLECUT ROWCOL 3 1 XPITCH 2 YPITCH 3 ;" ;
    
  LIBRARY LEF58_STACKVIARULE STRING "STACKVIARULE MY_VP5  VIA2_4X8_3X_USER VIA3_4X8_3X_USER VIA4_4X4_USER VIA5_4X4_USER VIA6_4X4_USER VIA7_4X4_USER VIA8_4X4_USER VIA9_3X4_USER VIA10_3X1_USER ;" ;      

  # Even heigher - up to this point we had 14 DRCs with only 3 on actuall M111-12 vias - BEST SO FAR
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA10_3X3_USER LAYER VIA10 CUTCLASS VSINGLECUT ROWCOL 3 3 XPITCH 2 YPITCH 3 ;" ;  
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA11_1X3_USER LAYER VIA11 CUTCLASS VSINGLECUT ROWCOL 1 3 XPITCH 4 YPITCH 3 MAXCELLEXTENSION 2 ;" ;  
    
  LIBRARY LEF58_STACKVIARULE STRING "STACKVIARULE MY_VP6  VIA2_4X8_3X_USER VIA3_4X8_3X_USER VIA4_4X4_USER VIA5_4X4_USER VIA6_4X4_USER VIA7_4X4_USER VIA8_4X4_USER VIA9_3X4_USER VIA10_3X3_USER VIA11_1X3_USER ;" ;      

  # Even heigher - up to this point we had 10 DRCs 
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA11_3X3_USER LAYER VIA11 CUTCLASS VSINGLECUT ROWCOL 3 3 XPITCH 6 YPITCH 3 MAXCELLEXTENSION 2 ;" ;    
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA12_3X1_USER LAYER VIA12 CUTCLASS VSINGLECUT ROWCOL 3 1 MAXCELLEXTENSION 2 ;" ;    
    
  LIBRARY LEF58_STACKVIARULE STRING "STACKVIARULE MY_VP7  VIA2_4X8_3X_USER VIA3_4X8_3X_USER VIA4_4X4_USER VIA5_4X4_USER VIA6_4X4_USER VIA7_4X4_USER VIA8_4X4_USER VIA9_3X4_USER VIA10_3X3_USER VIA11_3X3_USER VIA12_3X1_USER ;" ;        

  # Even heigher - Try to solve all the m11-m12 drcs
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA11_3X3_HP_USER LAYER VIA11 CUTCLASS VSINGLECUT ROWCOL 3 3 XPITCH 12 YPITCH 6 MAXCELLEXTENSION 2 ;" ;    
  LIBRARY LEF58_STACKVIALAYERRULE STRING "STACKVIALAYERRULE VIA12_3X1_HP_USER LAYER VIA12 CUTCLASS VSINGLECUT ROWCOL 3 1 XPITCH 12 YPITCH 6 MAXCELLEXTENSION 2 ;" ;    
    
  LIBRARY LEF58_STACKVIARULE STRING "STACKVIARULE MY_VP8  VIA2_4X8_3X_USER VIA3_4X8_3X_USER VIA4_4X4_USER VIA5_4X4_USER VIA6_4X4_USER VIA7_4X4_USER VIA8_4X4_USER VIA9_3X4_USER VIA10_3X3_USER VIA11_3X3_HP_USER VIA12_3X1_HP_USER ;" ;        
  

END PROPERTYDEFINITIONS


END LIBRARY
