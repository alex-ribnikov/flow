.SUBCKT rm1w p n
.ENDS

.SUBCKT rm2w p n
.ENDS
