SITE SPRBUF
    SIZE 27.132 BY 1.05 ;
    SYMMETRY Y ;
    CLASS CORE ;
END SPRBUF

SITE SPRBUF320R7
    SIZE 27.132 BY 9.24 ;
    SYMMETRY Y ;
    CLASS CORE ;
END SPRBUF320R7

SITE SPRBUF320T7
    SIZE 27.132 BY 1.47 ;
    SYMMETRY Y ;
    CLASS CORE ;
END SPRBUF320T7

SITE SPRBUF192R5
    SIZE 27.132 BY 5.88 ;
    SYMMETRY Y ;
    CLASS CORE ;
END SPRBUF192R5

SITE SPRBUF96R5
    SIZE 27.132 BY 3.36 ;
    SYMMETRY Y ;
    CLASS CORE ;
END SPRBUF96R5

SITE SPRBUF48G3
    SIZE 27.132 BY 0.63 ;
    SYMMETRY Y ;
    CLASS CORE ;
END SPRBUF48G3

SITE SPRBUF224R5
    SIZE 27.132 BY 6.72 ;
    SYMMETRY Y ;
    CLASS CORE ;
END SPRBUF224R5
